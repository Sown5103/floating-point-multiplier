module Sign_extend_R (In, Out);
input [47:0] In;
output [48:0] Out;
assign Out = In;
endmodule
